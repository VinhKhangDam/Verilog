module and_2 (
    input a ,b, 
    output result
);

and (result, a, b);
    
endmodule